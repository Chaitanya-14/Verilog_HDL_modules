module simple_and(f,a,b);
    input a,b;
    output f;
    assign f = a&b;
endmodule