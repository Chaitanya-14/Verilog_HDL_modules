`timescale 1ns / 1ns

module halfadder_tb;
    reg a,b;
    wire s,c;

    half_adder uut (.a(a),.b(b),.s(s),.c(c));

    initial
    begin
        $dumpfile("halfadder.vcd");
        $dumpvars(0,halfadder_tb);
        $monitor("Time=%0t|a=%b|b=%b|s=%b|c=%b",$time,a,b,s,c);
        a=0;b=0;#10;
        a=0;b=1;#10;
        a=1;b=0;#10;
        a=1;b=1;#10;
        $finish;
    end
endmodule

