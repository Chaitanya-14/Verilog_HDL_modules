module simple_not(f,a);
    input a;
    output f;
    assign f = ~a;
endmodule